`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:14:30 03/20/2015 
// Design Name: 
// Module Name:    UartReceiver 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module UartReceiver(
    input rxclk,
    input reset,
    input rxen,
    input rxin,
    input rxuld,
    output [7:0] rxrcvd
    );


endmodule
